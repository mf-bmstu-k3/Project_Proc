library verilog;
use verilog.vl_types.all;
entity CYY_AU_OP_with_RR_vlg_vec_tst is
end CYY_AU_OP_with_RR_vlg_vec_tst;
