library verilog;
use verilog.vl_types.all;
entity CYY_final_vlg_vec_tst is
end CYY_final_vlg_vec_tst;
